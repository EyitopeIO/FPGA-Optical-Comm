LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY rom IS
    PORT (
        data_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) ;  --32 bits
        addr: IN STD_LOGIC_VECTOR(8 DOWNTO 0)       --2^9 = 512
    );
END rom;

    --There are 404 elements

ARCHITECTURE romarch OF rom IS
    TYPE ro_memory IS ARRAY (0 TO 403) OF STD_LOGIC_VECTOR(31 DOWNTO 0) ;
    CONSTANT bytesel : ro_memory := (  

        x"7b7b224e",x"616d6522",x"3a226368",x"6576726f",x"6c657420",x"63686576",
        x"656c6c65",x"20636f6e",x"636f7572",x"73202873",x"7729222c",x"224d696c",
        x"65735f70",x"65725f47",x"616c6c6f",x"6e223a6e",x"756c6c2c",x"2243796c",
        x"696e6465",x"7273223a",x"382c2244",x"6973706c",x"6163656d",x"656e7422",
        x"3a333530",x"2c22486f",x"72736570",x"6f776572",x"223a3136",x"352c2257",
        x"65696768",x"745f696e",x"5f6c6273",x"223a3431",x"34322c22",x"41636365",
        x"6c657261",x"74696f6e",x"223a3131",x"2e352c22",x"59656172",x"223a2231",
        x"3937302d",x"30312d30",x"31222c22",x"4f726967",x"696e223a",x"22555341",
        x"227d2c7b",x"224e616d",x"65223a22",x"666f7264",x"20746f72",x"696e6f20",
        x"28737729",x"222c224d",x"696c6573",x"5f706572",x"5f47616c",x"6c6f6e22",
        x"3a6e756c",x"6c2c2243",x"796c696e",x"64657273",x"223a382c",x"22446973",
        x"706c6163",x"656d656e",x"74223a33",x"35312c22",x"486f7273",x"65706f77",
        x"6572223a",x"3135332c",x"22576569",x"6768745f",x"696e5f6c",x"6273223a",
        x"34303334",x"2c224163",x"63656c65",x"72617469",x"6f6e223a",x"31312c22",
        x"59656172",x"223a2231",x"3937302d",x"30312d30",x"31222c22",x"4f726967",
        x"696e223a",x"22555341",x"227d2c7b",x"224e616d",x"65223a22",x"616d6320",
        x"72656265",x"6c207373",x"74202873",x"7729222c",x"224d696c",x"65735f70",
        x"65725f47",x"616c6c6f",x"6e223a6e",x"756c6c2c",x"2243796c",x"696e6465",
        x"7273223a",x"382c2244",x"6973706c",x"6163656d",x"656e7422",x"3a333630",
        x"2c22486f",x"72736570",x"6f776572",x"223a3137",x"352c2257",x"65696768",
        x"745f696e",x"5f6c6273",x"223a3338",x"35302c22",x"41636365",x"6c657261",
        x"74696f6e",x"223a3131",x"2c225965",x"6172223a",x"22313937",x"302d3031",
        x"2d303122",x"2c224f72",x"6967696e",x"223a2255",x"5341227d",x"2c7b224e",
        x"616d6522",x"3a22646f",x"64676520",x"6368616c",x"6c656e67",x"65722073",
        x"65222c22",x"4d696c65",x"735f7065",x"725f4761",x"6c6c6f6e",x"223a3135",
        x"2c224379",x"6c696e64",x"65727322",x"3a382c22",x"44697370",x"6c616365",
        x"6d656e74",x"223a3338",x"332c2248",x"6f727365",x"706f7765",x"72223a31",
        x"37302c22",x"57656967",x"68745f69",x"6e5f6c62",x"73223a33",x"3536332c",
        x"22416363",x"656c6572",x"6174696f",x"6e223a31",x"302c2259",x"65617222",
        x"3a223139",x"37302d30",x"312d3031",x"222c224f",x"72696769",x"6e223a22",
        x"55534122",x"7d2c7b22",x"4e616d65",x"223a2270",x"6c796d6f",x"75746820",
        x"27637564",x"61203334",x"30222c22",x"4d696c65",x"735f7065",x"725f4761",
        x"6c6c6f6e",x"223a3134",x"2c224379",x"6c696e64",x"65727322",x"3a382c22",
        x"44697370",x"6c616365",x"6d656e74",x"223a3334",x"302c2248",x"6f727365",
        x"706f7765",x"72223a31",x"36302c22",x"57656967",x"68745f69",x"6e5f6c62",
        x"73223a33",x"3630392c",x"22416363",x"656c6572",x"6174696f",x"6e223a38",
        x"2c225965",x"6172223a",x"22313937",x"302d3031",x"2d303122",x"2c224f72",
        x"6967696e",x"223a2255",x"5341227d",x"2c7b224e",x"616d6522",x"3a22666f",
        x"7264206d",x"75737461",x"6e672062",x"6f737320",x"33303222",x"2c224d69",
        x"6c65735f",x"7065725f",x"47616c6c",x"6f6e223a",x"6e756c6c",x"2c224379",
        x"6c696e64",x"65727322",x"3a382c22",x"44697370",x"6c616365",x"6d656e74",
        x"223a3330",x"322c2248",x"6f727365",x"706f7765",x"72223a31",x"34302c22",
        x"57656967",x"68745f69",x"6e5f6c62",x"73223a33",x"3335332c",x"22416363",
        x"656c6572",x"6174696f",x"6e223a38",x"2c225965",x"6172223a",x"22313937",
        x"302d3031",x"2d303122",x"2c224f72",x"6967696e",x"223a2255",x"5341227d",
        x"2c7b224e",x"616d6522",x"3a226368",x"6576726f",x"6c657420",x"6d6f6e74",
        x"65206361",x"726c6f22",x"2c224d69",x"6c65735f",x"7065725f",x"47616c6c",
        x"6f6e223a",x"31352c22",x"43796c69",x"6e646572",x"73223a38",x"2c224469",
        x"73706c61",x"63656d65",x"6e74223a",x"3430302c",x"22486f72",x"7365706f",
        x"77657222",x"3a313530",x"2c225765",x"69676874",x"5f696e5f",x"6c627322",
        x"3a333736",x"312c2241",x"6363656c",x"65726174",x"696f6e22",x"3a392e35",
        x"2c225965",x"6172223a",x"22313937",x"302d3031",x"2d303122",x"2c224f72",
        x"6967696e",x"223a2255",x"5341227d",x"2c7b224e",x"616d6522",x"3a22746f",
        x"796f7461",x"20636f72",x"6f6e6120",x"6d61726b",x"20696922",x"2c224d69",
        x"6c65735f",x"7065725f",x"47616c6c",x"6f6e223a",x"32342c22",x"43796c69",
        x"6e646572",x"73223a34",x"2c224469",x"73706c61",x"63656d65",x"6e74223a",
        x"3131332c",x"22486f72",x"7365706f",x"77657222",x"3a39352c",x"22576569",
        x"6768745f",x"696e5f6c",x"6273223a",x"32333732",x"2c224163",x"63656c65",
        x"72617469",x"6f6e223a",x"31352c22",x"59656172",x"223a2231",x"3937302d",
        x"30312d30",x"31222c22",x"4f726967",x"696e223a",x"224a6170",x"616e227d",
        x"2c7b224e",x"616d6522",x"3a22706c",x"796d6f75",x"74682064",x"75737465",
        x"72222c22",x"4d696c65",x"735f7065",x"725f4761",x"6c6c6f6e",x"223a3232",
        x"2c224379",x"6c696e64",x"65727322",x"3a362c22",x"44697370",x"6c616365",
        x"6d656e74",x"223a3139",x"382c2248",x"6f727365",x"706f7765",x"72223a39",
        x"352c2257",x"65696768",x"745f696e",x"5f6c6273",x"223a3238",x"33332c22",
        x"41636365",x"6c657261",x"74696f6e",x"223a3135",x"2e352c22",x"59656172",
        x"223a2231",x"3937302d",x"30312d30",x"31222c22",x"4f726967",x"696e223a",
        x"22555341",x"ffffffff"
    );
BEGIN
    data_out <= bytesel(TO_INTEGER(UNSIGNED(addr))) WHEN UNSIGNED(addr) < 404 ELSE x"FFFFFFFF" ;
END romarch ;
                            

